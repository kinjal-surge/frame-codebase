component osc_ip is
    port(
        hf_out_en_i: in std_logic;
        hf_clk_out_o: out std_logic
    );
end component;

__: osc_ip port map(
    hf_out_en_i=>,
    hf_clk_out_o=>
);
